module picture_gen #(parameter WIDTH=8) (
    input logic [3:0] id,
    output logic [7:0][WIDTH-1:0] pic 
);
    always_comb begin
        case (id) 
            4'd0 : begin
                pic = {
                    8'b00111100, 
                    8'b01100110,
                    8'b01100110,
                    8'b01100110,
                    8'b01100110,
                    8'b01100110,
                    8'b00111100,
                    8'b00000000
                };
            end
            4'd1 : begin
                pic = {
                    8'b00011000,
                    8'b00111000,
                    8'b00011000,
                    8'b00011000,
                    8'b00011000,
                    8'b00011000,
                    8'b00111100,
                    8'b00000000
                };
            end
            4'd2 : begin
                pic = {
                    8'b00111100,
                    8'b01100110,
                    8'b00000110,
                    8'b00011100,
                    8'b00110000,
                    8'b01100000,
                    8'b01111110,
                    8'b00000000
                };
            end
            4'd3 : begin
                pic = {
                    8'b00111100,
                    8'b01100110,
                    8'b00000110,
                    8'b00011100,
                    8'b00000110,
                    8'b01100110,
                    8'b00111100,
                    8'b00000000
                };
            end
            4'd4 : begin
                pic = {
                    8'b01100110,
                    8'b01100110,
                    8'b01100110,
                    8'b01111110,
                    8'b00000110,
                    8'b00000110,
                    8'b00000110,
                    8'b00000000
                };
            end
            4'd5 : begin
                pic = {
                    8'b01111110,
                    8'b01100000,
                    8'b01111100,
                    8'b00000110,
                    8'b00000110,
                    8'b01100110,
                    8'b00111100,
                    8'b00000000
                };
            end
            4'd6 : begin
                pic = {
                    8'b00111100,
                    8'b01100110,
                    8'b01100000,
                    8'b01111100,
                    8'b01100110,
                    8'b01100110,
                    8'b00111100,
                    8'b00000000
                };
            end
            4'd7 : begin
                pic = {
                    8'b01111110,
                    8'b00000110,
                    8'b00001100,
                    8'b00011000,
                    8'b00011000,
                    8'b00011000,
                    8'b00011000,
                    8'b00000000
                };
            end
            4'd8 : begin // cat
                 pic = {
                    8'b01000010,
                    8'b10100101,
                    8'b10011001,
                    8'b01111110,
                    8'b10000001,
                    8'b10100101,
                    8'b10000001,
                    8'b01111110
                };
            end
            4'd9 : begin // WIN
                 pic = {
                    16'b1000101110100010,
                    16'b1000100100110010,
                    16'b1000100100101010,
                    16'b1010100100100110,
                    16'b0101001110100010,
                    16'd0,
                    16'd0,
                    16'd0
                };
            end
            default : begin
                pic = {
                    8'b01111110,
                    8'b01111110,
                    8'b01111110,
                    8'b01111110,
                    8'b01111110,
                    8'b01111110,
                    8'b01111110,
                    8'b01111110
                };
            end
        endcase
    end
endmodule